module myXOR(input x,y, output z);   //kendi modulümüzü oluşturduk.

	xor x1(z,x,y);
	
endmodule	
