module example(A,B,C,Z);


		input A,B,C;
		output Z;

		and a1(Z,A,B,C);
	
endmodule 