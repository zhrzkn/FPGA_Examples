module trial(
   input [4:0] IN,
   input in1,in2,in3,in4,
	output [4:0] OUT,
	output o1,o2);
	
endmodule	